library ieee;
library work;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.ALL;
use IEEE.STD_LOGIC_TEXTIO.all;
use STD.TEXTIO.all;
use work.opcodes.all;
--use work.Components.all;


entity dft is
		generic(ROWS  : 	integer := 15;
				COLUMNS :   integer := 3);
		port(	);
end entity;


architecture arch of fft_dfg is





end arch;